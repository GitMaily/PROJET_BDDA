�� sr Catalog05�1��S I compteurRelationL listRIt Ljava/util/ArrayList;L patht Ljava/lang/String;xp    sr java.util.ArrayListx����a� I sizexp   w   sr RelationInfo�W����e I nb_colL headert LPageId;L headerPageIdq ~ L nomq ~ L nom_colq ~ xp   psr PageId�!��K� I FileIdxI PageIdxxp        t Profssq ~    w   sr ColInfov���Y�W L nom_colq ~ L type_colq ~ xpt NOMt VARCHAR(10)sq ~ t UEq ~ xsq ~    pq ~ 
t 	Etudiantssq ~    w   sq ~ q ~ q ~ sq ~ t PRENOMq ~ xxt _C:\Users\milly\Desktop\PROJET_BDDA\PROJET_BDDA_LAVALLEE_TANGUY_CIAVALDINI_MARZOUK\DB\catalog.sv