�� {sr  java.io.NotSerializableException(Vx �5  xr java.io.ObjectStreamExceptiond��k�9��  xr java.io.IOExceptionl�sde%�  xr java.lang.Exception��>;�  xr java.lang.Throwable��5'9w�� L causet Ljava/lang/Throwable;L detailMessaget Ljava/lang/String;[ 
stackTracet [Ljava/lang/StackTraceElement;L suppressedExceptionst Ljava/util/List;xpq ~ 	t Catalogur [Ljava.lang.StackTraceElement;F*<<�"9  xp   sr java.lang.StackTraceElementa	Ś&6݅ B formatI 
lineNumberL classLoaderNameq ~ L declaringClassq ~ L fileNameq ~ L 
methodNameq ~ L 
moduleNameq ~ L moduleVersionq ~ xp  �pt java.io.ObjectOutputStreamt ObjectOutputStream.javat writeObject0t 	java.baset 17.0.4.1sq ~   ^pq ~ q ~ t writeObjectq ~ q ~ sq ~    (t appq ~ 
t Catalog.javat Finishppsq ~    
q ~ t TestCatalogt TestCatalog.javat addRelationTestppsq ~    q ~ q ~ q ~ t mainppsr java.util.Collections$EmptyListz��<���  xpx