�� sr Catalog05�1��S I compteurRelationL listRIt Ljava/util/ArrayList;L patht Ljava/lang/String;xp    sr java.util.ArrayListx����a� I sizexp   w   sr RelationInfo�W����e I nb_colL headert LPageId;L headerPageIdq ~ L nomq ~ L nom_colq ~ xp   psr PageId�!��K� I FileIdxI PageIdxxp        t Ssq ~    w   sr ColInfov���Y�W L nom_colq ~ L type_colq ~ xpt C1t INTEGERsq ~ t C2t REALsq ~ t C3t INTEGERsq ~ t C4t INTEGERsq ~ t C5t INTEGERxxt eC:\\Users\\milly\\Desktop\\PROJET_BDDA\\PROJET_BDDA_LAVALLEE_TANGUY_CIAVALDINI_MARZOUK\\DB\catalog.sv