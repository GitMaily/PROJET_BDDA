�� sr Catalog05�1��S I compteurRelationL listRIt Ljava/util/ArrayList;L patht Ljava/lang/String;xp    sr java.util.ArrayListx����a� I sizexp    w    xt _C:\Users\milly\Desktop\PROJET_BDDA\PROJET_BDDA_LAVALLEE_TANGUY_CIAVALDINI_MARZOUK\DB\catalog.sv